//  1 bit ALU
module ALU_1(A, B, C_in, cntrl, C_out, S);

	input logic A, B, C_in;
	input logic [2:0] cntrl;
	output logic C_out, S;

endmodule
