`timescale 1ns/10ps

// 64 bit or
module or_64();


endmodule