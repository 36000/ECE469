`timescale 1ns/10ps

//  input flags, output conditional signals
module ();

endmodule